//Instructions
`DEFINE LD     6'b011000
`DEFINE ST     6'b011001
`DEFINE JMP    6'b011011
`DEFINE BEQ    6'b011100
`DEFINE BNE    6'b011101
`DEFINE LDR    6'b011111
`DEFINE ADD    6'b100000
`DEFINE SUB    6'b100001
`DEFINE MUL    6'b100010
`DEFINE DIV    6'b100011
`DEFINE CMPEQ  6'b100100
`DEFINE CMPLT  6'b100101
`DEFINE CMPLE  6'b100110
`DEFINE AND    6'b101000
`DEFINE OR     6'b101001
`DEFINE XOR    6'b101010
`DEFINE XNOR   6'b101011
`DEFINE SHL    6'b101100
`DEFINE SHR    6'b101101
`DEFINE SRA    6'b101110
`DEFINE ADDC   6'b101000
`DEFINE SUBC   6'b110001
`DEFINE MULC   6'b110010
`DEFINE DIVC   6'b110011
`DEFINE CMPEQC 6'b110100
`DEFINE CMPLTC 6'b110101
`DEFINE CMPLEC 6'b110110
`DEFINE ANDC   6'b111000
`DEFINE ORC    6'b111001
`DEFINE XORC   6'b111010
`DEFINE XNORC  6'b111011
`DEFINE SHLC   6'b111100
`DEFINE SHRC   6'b111101
`DEFINE SRAC   6'b111110
