//Instructions
`define LD     6'b011000
`define ST     6'b011001
`define DISP   6'b011010
`define JMP    6'b011011
`define BEQ    6'b011100
`define BNE    6'b011101
`define DISPC  6'b011110
`define LDR    6'b011111
`define ADD    6'b100000
`define SUB    6'b100001
`define MUL    6'b100010
`define DIV    6'b100011
`define CMPEQ  6'b100100
`define CMPLT  6'b100101
`define CMPLE  6'b100110
`define AND    6'b101000
`define OR     6'b101001
`define XOR    6'b101010
`define XNOR   6'b101011
`define SHL    6'b101100
`define SHR    6'b101101
`define SRA    6'b101110
`define ADDC   6'b101000
`define SUBC   6'b110001
`define MULC   6'b110010
`define DIVC   6'b110011
`define CMPEQC 6'b110100
`define CMPLTC 6'b110101
`define CMPLEC 6'b110110
`define ANDC   6'b111000
`define ORC    6'b111001
`define XORC   6'b111010
`define XNORC  6'b111011
`define SHLC   6'b111100
`define SHRC   6'b111101
`define SRAC   6'b111110
