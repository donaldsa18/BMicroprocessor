`DEFINE DWIDTH 32
`DEFINE MEMDEPTH 1024
`DEFINE AWIDTH $clog2(MEMDEPTH)
`DEFINE CPUAWIDTH 16
`DEFINE NUM_REGS 32