parameter DWIDTH = 32;
parameter MEMDEPTH = 1024;
parameter AWIDTH = $clog2(MEMDEPTH);
parameter CPUAWIDTH = 16;
parameter NUM_REGS = 32;